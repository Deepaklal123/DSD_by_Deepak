`timescale 1ns / 1ps

module And_Gate(input a,b, output c );

and and1 (c, a,b);
endmodule
